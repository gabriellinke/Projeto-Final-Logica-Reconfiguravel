-- system_0_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2023.06.24.22:14:45

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_0_tb is
end entity system_0_tb;

architecture rtl of system_0_tb is
	component system_0 is
		port (
			clk_50                               : in    std_logic                     := 'X';             -- clk
			bidir_port_to_and_from_the_SD_DAT    : inout std_logic                     := 'X';             -- export
			out_port_from_the_led_red            : out   std_logic_vector(17 downto 0);                    -- export
			zs_addr_from_the_sdram_0             : out   std_logic_vector(11 downto 0);                    -- addr
			zs_ba_from_the_sdram_0               : out   std_logic_vector(1 downto 0);                     -- ba
			zs_cas_n_from_the_sdram_0            : out   std_logic;                                        -- cas_n
			zs_cke_from_the_sdram_0              : out   std_logic;                                        -- cke
			zs_cs_n_from_the_sdram_0             : out   std_logic;                                        -- cs_n
			zs_dq_to_and_from_the_sdram_0        : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			zs_dqm_from_the_sdram_0              : out   std_logic_vector(1 downto 0);                     -- dqm
			zs_ras_n_from_the_sdram_0            : out   std_logic;                                        -- ras_n
			zs_we_n_from_the_sdram_0             : out   std_logic;                                        -- we_n
			tri_state_bridge_0_data              : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			tri_state_bridge_0_readn             : out   std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0           : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address           : out   std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0          : out   std_logic_vector(0 downto 0);                     -- select_n_to_the_cfi_flash_0
			reset_n                              : in    std_logic                     := 'X';             -- reset_n
			bidir_port_to_and_from_the_SD_CMD    : inout std_logic                     := 'X';             -- export
			in_port_to_the_button_pio            : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			USB_DATA_to_and_from_the_ISP1362     : inout std_logic_vector(15 downto 0) := (others => 'X'); -- DATA
			USB_ADDR_from_the_ISP1362            : out   std_logic_vector(1 downto 0);                     -- ADDR
			USB_RD_N_from_the_ISP1362            : out   std_logic;                                        -- RD_N
			USB_WR_N_from_the_ISP1362            : out   std_logic;                                        -- WR_N
			USB_CS_N_from_the_ISP1362            : out   std_logic;                                        -- CS_N
			USB_RST_N_from_the_ISP1362           : out   std_logic;                                        -- RST_N
			USB_INT0_to_the_ISP1362              : in    std_logic                     := 'X';             -- INT0
			USB_INT1_to_the_ISP1362              : in    std_logic                     := 'X';             -- INT1
			out_port_from_the_SD_CLK             : out   std_logic;                                        -- export
			out_port_from_the_led_green          : out   std_logic_vector(8 downto 0);                     -- export
			in_port_to_the_switch_pio            : in    std_logic_vector(17 downto 0) := (others => 'X'); -- export
			LCD_RS_from_the_lcd_16207_0          : out   std_logic;                                        -- RS
			LCD_RW_from_the_lcd_16207_0          : out   std_logic;                                        -- RW
			LCD_data_to_and_from_the_lcd_16207_0 : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			LCD_E_from_the_lcd_16207_0           : out   std_logic;                                        -- E
			rxd_to_the_uart_0                    : in    std_logic                     := 'X';             -- rxd
			txd_from_the_uart_0                  : out   std_logic;                                        -- txd
			audio_0_oAUD_DATA                    : out   std_logic;                                        -- oAUD_DATA
			audio_0_oAUD_LRCK                    : out   std_logic;                                        -- oAUD_LRCK
			audio_0_oAUD_BCK                     : out   std_logic;                                        -- oAUD_BCK
			audio_0_oAUD_XCK                     : out   std_logic;                                        -- oAUD_XCK
			audio_0_iCLK_18_4                    : in    std_logic                     := 'X';             -- iCLK_18_4
			vga_0_VGA_R                          : out   std_logic_vector(9 downto 0);                     -- VGA_R
			vga_0_VGA_G                          : out   std_logic_vector(9 downto 0);                     -- VGA_G
			vga_0_VGA_B                          : out   std_logic_vector(9 downto 0);                     -- VGA_B
			vga_0_VGA_HS                         : out   std_logic;                                        -- VGA_HS
			vga_0_VGA_VS                         : out   std_logic;                                        -- VGA_VS
			vga_0_VGA_SYNC                       : out   std_logic;                                        -- VGA_SYNC
			vga_0_VGA_BLANK                      : out   std_logic;                                        -- VGA_BLANK
			vga_0_VGA_CLK                        : out   std_logic;                                        -- VGA_CLK
			vga_0_iCLK_25                        : in    std_logic                     := 'X';             -- iCLK_25
			dm9000a_iOSC_50                      : in    std_logic                     := 'X';             -- iOSC_50
			dm9000a_ENET_DATA                    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- ENET_DATA
			dm9000a_ENET_CMD                     : out   std_logic;                                        -- ENET_CMD
			dm9000a_ENET_RD_N                    : out   std_logic;                                        -- ENET_RD_N
			dm9000a_ENET_WR_N                    : out   std_logic;                                        -- ENET_WR_N
			dm9000a_ENET_CS_N                    : out   std_logic;                                        -- ENET_CS_N
			dm9000a_ENET_RST_N                   : out   std_logic;                                        -- ENET_RST_N
			dm9000a_ENET_CLK                     : out   std_logic;                                        -- ENET_CLK
			dm9000a_ENET_INT                     : in    std_logic                     := 'X';             -- ENET_INT
			seg7_display_oSEG0                   : out   std_logic_vector(6 downto 0);                     -- oSEG0
			seg7_display_oSEG1                   : out   std_logic_vector(6 downto 0);                     -- oSEG1
			seg7_display_oSEG2                   : out   std_logic_vector(6 downto 0);                     -- oSEG2
			seg7_display_oSEG3                   : out   std_logic_vector(6 downto 0);                     -- oSEG3
			seg7_display_oSEG4                   : out   std_logic_vector(6 downto 0);                     -- oSEG4
			seg7_display_oSEG5                   : out   std_logic_vector(6 downto 0);                     -- oSEG5
			seg7_display_oSEG6                   : out   std_logic_vector(6 downto 0);                     -- oSEG6
			seg7_display_oSEG7                   : out   std_logic_vector(6 downto 0)                      -- oSEG7
		);
	end component system_0;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_export : inout std_logic := 'X'  -- export
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : in std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_export : out std_logic_vector(3 downto 0)   -- export
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_DATA  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- DATA
			sig_ADDR  : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ADDR
			sig_RD_N  : in    std_logic                     := 'X';             -- RD_N
			sig_WR_N  : in    std_logic                     := 'X';             -- WR_N
			sig_CS_N  : in    std_logic                     := 'X';             -- CS_N
			sig_RST_N : in    std_logic                     := 'X';             -- RST_N
			sig_INT0  : out   std_logic;                                        -- INT0
			sig_INT1  : out   std_logic                                         -- INT1
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_export : in std_logic := 'X'  -- export
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			sig_export : in std_logic_vector(8 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0006;

	component altera_conduit_bfm_0007 is
		port (
			sig_export : out std_logic_vector(17 downto 0)   -- export
		);
	end component altera_conduit_bfm_0007;

	component altera_conduit_bfm_0008 is
		port (
			sig_RS   : in    std_logic                    := 'X';             -- RS
			sig_RW   : in    std_logic                    := 'X';             -- RW
			sig_data : inout std_logic_vector(7 downto 0) := (others => 'X'); -- data
			sig_E    : in    std_logic                    := 'X'              -- E
		);
	end component altera_conduit_bfm_0008;

	component altera_conduit_bfm_0009 is
		port (
			sig_rxd : out std_logic;        -- rxd
			sig_txd : in  std_logic := 'X'  -- txd
		);
	end component altera_conduit_bfm_0009;

	component altera_conduit_bfm_0010 is
		port (
			sig_oAUD_DATA : in  std_logic := 'X'; -- oAUD_DATA
			sig_oAUD_LRCK : in  std_logic := 'X'; -- oAUD_LRCK
			sig_oAUD_BCK  : in  std_logic := 'X'; -- oAUD_BCK
			sig_oAUD_XCK  : in  std_logic := 'X'; -- oAUD_XCK
			sig_iCLK_18_4 : out std_logic         -- iCLK_18_4
		);
	end component altera_conduit_bfm_0010;

	component altera_conduit_bfm_0011 is
		port (
			sig_VGA_R     : in  std_logic_vector(9 downto 0) := (others => 'X'); -- VGA_R
			sig_VGA_G     : in  std_logic_vector(9 downto 0) := (others => 'X'); -- VGA_G
			sig_VGA_B     : in  std_logic_vector(9 downto 0) := (others => 'X'); -- VGA_B
			sig_VGA_HS    : in  std_logic                    := 'X';             -- VGA_HS
			sig_VGA_VS    : in  std_logic                    := 'X';             -- VGA_VS
			sig_VGA_SYNC  : in  std_logic                    := 'X';             -- VGA_SYNC
			sig_VGA_BLANK : in  std_logic                    := 'X';             -- VGA_BLANK
			sig_VGA_CLK   : in  std_logic                    := 'X';             -- VGA_CLK
			sig_iCLK_25   : out std_logic                                        -- iCLK_25
		);
	end component altera_conduit_bfm_0011;

	component altera_conduit_bfm_0012 is
		port (
			sig_iOSC_50    : out   std_logic;                                        -- iOSC_50
			sig_ENET_DATA  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- ENET_DATA
			sig_ENET_CMD   : in    std_logic                     := 'X';             -- ENET_CMD
			sig_ENET_RD_N  : in    std_logic                     := 'X';             -- ENET_RD_N
			sig_ENET_WR_N  : in    std_logic                     := 'X';             -- ENET_WR_N
			sig_ENET_CS_N  : in    std_logic                     := 'X';             -- ENET_CS_N
			sig_ENET_RST_N : in    std_logic                     := 'X';             -- ENET_RST_N
			sig_ENET_CLK   : in    std_logic                     := 'X';             -- ENET_CLK
			sig_ENET_INT   : out   std_logic                                         -- ENET_INT
		);
	end component altera_conduit_bfm_0012;

	component altera_conduit_bfm_0013 is
		port (
			sig_oSEG0 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG0
			sig_oSEG1 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG1
			sig_oSEG2 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG2
			sig_oSEG3 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG3
			sig_oSEG4 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG4
			sig_oSEG5 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG5
			sig_oSEG6 : in std_logic_vector(6 downto 0) := (others => 'X'); -- oSEG6
			sig_oSEG7 : in std_logic_vector(6 downto 0) := (others => 'X')  -- oSEG7
		);
	end component altera_conduit_bfm_0013;

	component altera_sdram_partner_module is
		port (
			clk      : in    std_logic                     := 'X';             -- clk
			zs_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			zs_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			zs_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			zs_cas_n : in    std_logic                     := 'X';             -- cas_n
			zs_cke   : in    std_logic                     := 'X';             -- cke
			zs_cs_n  : in    std_logic                     := 'X';             -- cs_n
			zs_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			zs_ras_n : in    std_logic                     := 'X';             -- ras_n
			zs_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_sdram_partner_module;

	component altera_tristate_conduit_bridge_translator is
		port (
			in_tri_state_bridge_0_data     : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			in_tri_state_bridge_0_readn    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_address  : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tri_state_bridge_0_address
			in_select_n_to_the_cfi_flash_0 : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_0
			tri_state_bridge_0_data        : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			tri_state_bridge_0_readn       : out   std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0     : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address     : out   std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0    : out   std_logic_vector(0 downto 0)                      -- select_n_to_the_cfi_flash_0
		);
	end component altera_tristate_conduit_bridge_translator;

	component altera_conduit_pin_divider is
		port (
			in_tri_state_bridge_0_address    : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tri_state_bridge_0_address
			in_tri_state_bridge_0_readn      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_data       : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			in_select_n_to_the_cfi_flash_0   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_0
			cfi_flash_0_tcm_address_out      : out   std_logic_vector(21 downto 0);                    -- tcm_address_out
			cfi_flash_0_tcm_read_n_out       : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			cfi_flash_0_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			cfi_flash_0_tcm_data_out         : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tcm_data_out
			cfi_flash_0_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component altera_conduit_pin_divider;

	component altera_external_memory_bfm_vhdl is
		generic (
			USE_CHIPSELECT           : integer := 1;
			USE_WRITE                : integer := 1;
			USE_READ                 : integer := 1;
			USE_OUTPUTENABLE         : integer := 1;
			USE_BEGINTRANSFER        : integer := 1;
			ACTIVE_LOW_BYTEENABLE    : integer := 0;
			ACTIVE_LOW_CHIPSELECT    : integer := 0;
			ACTIVE_LOW_WRITE         : integer := 0;
			ACTIVE_LOW_READ          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE  : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER : integer := 0;
			ACTIVE_LOW_RESET         : integer := 0;
			CDT_ADDRESS_W            : integer := 8;
			CDT_SYMBOL_W             : integer := 8;
			CDT_NUMSYMBOLS           : integer := 4;
			INIT_FILE                : string  := "altera_external_memory_bfm.hex";
			CDT_READ_LATENCY         : integer := 0;
			VHDL_ID                  : integer := 0
		);
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			cdt_write         : in    std_logic                     := 'X';             -- tcm_write_n_out
			cdt_read          : in    std_logic                     := 'X';             -- tcm_read_n_out
			cdt_chipselect    : in    std_logic                     := 'X';             -- tcm_chipselect_n_out
			cdt_address       : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tcm_address_out
			cdt_data_io       : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tcm_data_out
			cdt_outputenable  : in    std_logic                     := 'X';             -- tcm_outputenable_out
			cdt_begintransfer : in    std_logic                     := 'X';             -- tcm_begintransfer_out
			cdt_byteenable    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_byteenable_out
			cdt_reset         : in    std_logic                     := 'X'              -- tcm_reset_out
		);
	end component altera_external_memory_bfm_vhdl;

	signal system_0_inst_clk_50_clk_in_bfm_clk_clk                                         : std_logic;                     -- system_0_inst_clk_50_clk_in_bfm:clk -> [cfi_flash_0_external_mem_bfm:clk, sdram_0_my_partner:clk, system_0_inst:clk_50, system_0_inst_merged_resets_in_reset_bfm:clk]
	signal system_0_inst_merged_resets_in_reset_bfm_reset_reset                            : std_logic;                     -- system_0_inst_merged_resets_in_reset_bfm:reset -> system_0_inst:reset_n
	signal system_0_inst_sd_dat_external_connection_export                                 : std_logic;                     -- [] -> [system_0_inst:bidir_port_to_and_from_the_SD_DAT, system_0_inst_SD_DAT_external_connection_bfm:sig_export]
	signal system_0_inst_led_red_external_connection_export                                : std_logic_vector(17 downto 0); -- system_0_inst:out_port_from_the_led_red -> system_0_inst_led_red_external_connection_bfm:sig_export
	signal system_0_inst_sd_cmd_external_connection_export                                 : std_logic;                     -- [] -> [system_0_inst:bidir_port_to_and_from_the_SD_CMD, system_0_inst_SD_CMD_external_connection_bfm:sig_export]
	signal system_0_inst_button_pio_external_connection_bfm_conduit_export                 : std_logic_vector(3 downto 0);  -- system_0_inst_button_pio_external_connection_bfm:sig_export -> system_0_inst:in_port_to_the_button_pio
	signal system_0_inst_isp1362_conduit_end_wr_n                                          : std_logic;                     -- system_0_inst:USB_WR_N_from_the_ISP1362 -> system_0_inst_ISP1362_conduit_end_bfm:sig_WR_N
	signal system_0_inst_isp1362_conduit_end_bfm_conduit_int0                              : std_logic;                     -- system_0_inst_ISP1362_conduit_end_bfm:sig_INT0 -> system_0_inst:USB_INT0_to_the_ISP1362
	signal system_0_inst_isp1362_conduit_end_cs_n                                          : std_logic;                     -- system_0_inst:USB_CS_N_from_the_ISP1362 -> system_0_inst_ISP1362_conduit_end_bfm:sig_CS_N
	signal system_0_inst_isp1362_conduit_end_bfm_conduit_int1                              : std_logic;                     -- system_0_inst_ISP1362_conduit_end_bfm:sig_INT1 -> system_0_inst:USB_INT1_to_the_ISP1362
	signal system_0_inst_isp1362_conduit_end_addr                                          : std_logic_vector(1 downto 0);  -- system_0_inst:USB_ADDR_from_the_ISP1362 -> system_0_inst_ISP1362_conduit_end_bfm:sig_ADDR
	signal system_0_inst_isp1362_conduit_end_data                                          : std_logic_vector(15 downto 0); -- [] -> [system_0_inst:USB_DATA_to_and_from_the_ISP1362, system_0_inst_ISP1362_conduit_end_bfm:sig_DATA]
	signal system_0_inst_isp1362_conduit_end_rst_n                                         : std_logic;                     -- system_0_inst:USB_RST_N_from_the_ISP1362 -> system_0_inst_ISP1362_conduit_end_bfm:sig_RST_N
	signal system_0_inst_isp1362_conduit_end_rd_n                                          : std_logic;                     -- system_0_inst:USB_RD_N_from_the_ISP1362 -> system_0_inst_ISP1362_conduit_end_bfm:sig_RD_N
	signal system_0_inst_sd_clk_external_connection_export                                 : std_logic;                     -- system_0_inst:out_port_from_the_SD_CLK -> system_0_inst_SD_CLK_external_connection_bfm:sig_export
	signal system_0_inst_led_green_external_connection_export                              : std_logic_vector(8 downto 0);  -- system_0_inst:out_port_from_the_led_green -> system_0_inst_led_green_external_connection_bfm:sig_export
	signal system_0_inst_switch_pio_external_connection_bfm_conduit_export                 : std_logic_vector(17 downto 0); -- system_0_inst_switch_pio_external_connection_bfm:sig_export -> system_0_inst:in_port_to_the_switch_pio
	signal system_0_inst_lcd_16207_0_external_e                                            : std_logic;                     -- system_0_inst:LCD_E_from_the_lcd_16207_0 -> system_0_inst_lcd_16207_0_external_bfm:sig_E
	signal system_0_inst_lcd_16207_0_external_rs                                           : std_logic;                     -- system_0_inst:LCD_RS_from_the_lcd_16207_0 -> system_0_inst_lcd_16207_0_external_bfm:sig_RS
	signal system_0_inst_lcd_16207_0_external_rw                                           : std_logic;                     -- system_0_inst:LCD_RW_from_the_lcd_16207_0 -> system_0_inst_lcd_16207_0_external_bfm:sig_RW
	signal system_0_inst_lcd_16207_0_external_data                                         : std_logic_vector(7 downto 0);  -- [] -> [system_0_inst:LCD_data_to_and_from_the_lcd_16207_0, system_0_inst_lcd_16207_0_external_bfm:sig_data]
	signal system_0_inst_uart_0_external_connection_bfm_conduit_rxd                        : std_logic;                     -- system_0_inst_uart_0_external_connection_bfm:sig_rxd -> system_0_inst:rxd_to_the_uart_0
	signal system_0_inst_uart_0_external_connection_txd                                    : std_logic;                     -- system_0_inst:txd_from_the_uart_0 -> system_0_inst_uart_0_external_connection_bfm:sig_txd
	signal system_0_inst_audio_0_oaud_data                                                 : std_logic;                     -- system_0_inst:audio_0_oAUD_DATA -> system_0_inst_audio_0_bfm:sig_oAUD_DATA
	signal system_0_inst_audio_0_oaud_lrck                                                 : std_logic;                     -- system_0_inst:audio_0_oAUD_LRCK -> system_0_inst_audio_0_bfm:sig_oAUD_LRCK
	signal system_0_inst_audio_0_bfm_conduit_iclk_18_4                                     : std_logic;                     -- system_0_inst_audio_0_bfm:sig_iCLK_18_4 -> system_0_inst:audio_0_iCLK_18_4
	signal system_0_inst_audio_0_oaud_bck                                                  : std_logic;                     -- system_0_inst:audio_0_oAUD_BCK -> system_0_inst_audio_0_bfm:sig_oAUD_BCK
	signal system_0_inst_audio_0_oaud_xck                                                  : std_logic;                     -- system_0_inst:audio_0_oAUD_XCK -> system_0_inst_audio_0_bfm:sig_oAUD_XCK
	signal system_0_inst_vga_0_vga_vs                                                      : std_logic;                     -- system_0_inst:vga_0_VGA_VS -> system_0_inst_vga_0_bfm:sig_VGA_VS
	signal system_0_inst_vga_0_vga_r                                                       : std_logic_vector(9 downto 0);  -- system_0_inst:vga_0_VGA_R -> system_0_inst_vga_0_bfm:sig_VGA_R
	signal system_0_inst_vga_0_vga_g                                                       : std_logic_vector(9 downto 0);  -- system_0_inst:vga_0_VGA_G -> system_0_inst_vga_0_bfm:sig_VGA_G
	signal system_0_inst_vga_0_vga_sync                                                    : std_logic;                     -- system_0_inst:vga_0_VGA_SYNC -> system_0_inst_vga_0_bfm:sig_VGA_SYNC
	signal system_0_inst_vga_0_vga_clk                                                     : std_logic;                     -- system_0_inst:vga_0_VGA_CLK -> system_0_inst_vga_0_bfm:sig_VGA_CLK
	signal system_0_inst_vga_0_vga_blank                                                   : std_logic;                     -- system_0_inst:vga_0_VGA_BLANK -> system_0_inst_vga_0_bfm:sig_VGA_BLANK
	signal system_0_inst_vga_0_bfm_conduit_iclk_25                                         : std_logic;                     -- system_0_inst_vga_0_bfm:sig_iCLK_25 -> system_0_inst:vga_0_iCLK_25
	signal system_0_inst_vga_0_vga_hs                                                      : std_logic;                     -- system_0_inst:vga_0_VGA_HS -> system_0_inst_vga_0_bfm:sig_VGA_HS
	signal system_0_inst_vga_0_vga_b                                                       : std_logic_vector(9 downto 0);  -- system_0_inst:vga_0_VGA_B -> system_0_inst_vga_0_bfm:sig_VGA_B
	signal system_0_inst_dm9000a_enet_rd_n                                                 : std_logic;                     -- system_0_inst:dm9000a_ENET_RD_N -> system_0_inst_dm9000a_bfm:sig_ENET_RD_N
	signal system_0_inst_dm9000a_enet_wr_n                                                 : std_logic;                     -- system_0_inst:dm9000a_ENET_WR_N -> system_0_inst_dm9000a_bfm:sig_ENET_WR_N
	signal system_0_inst_dm9000a_enet_cmd                                                  : std_logic;                     -- system_0_inst:dm9000a_ENET_CMD -> system_0_inst_dm9000a_bfm:sig_ENET_CMD
	signal system_0_inst_dm9000a_bfm_conduit_enet_int                                      : std_logic;                     -- system_0_inst_dm9000a_bfm:sig_ENET_INT -> system_0_inst:dm9000a_ENET_INT
	signal system_0_inst_dm9000a_enet_cs_n                                                 : std_logic;                     -- system_0_inst:dm9000a_ENET_CS_N -> system_0_inst_dm9000a_bfm:sig_ENET_CS_N
	signal system_0_inst_dm9000a_bfm_conduit_iosc_50                                       : std_logic;                     -- system_0_inst_dm9000a_bfm:sig_iOSC_50 -> system_0_inst:dm9000a_iOSC_50
	signal system_0_inst_dm9000a_enet_rst_n                                                : std_logic;                     -- system_0_inst:dm9000a_ENET_RST_N -> system_0_inst_dm9000a_bfm:sig_ENET_RST_N
	signal system_0_inst_dm9000a_enet_clk                                                  : std_logic;                     -- system_0_inst:dm9000a_ENET_CLK -> system_0_inst_dm9000a_bfm:sig_ENET_CLK
	signal system_0_inst_dm9000a_enet_data                                                 : std_logic_vector(15 downto 0); -- [] -> [system_0_inst:dm9000a_ENET_DATA, system_0_inst_dm9000a_bfm:sig_ENET_DATA]
	signal system_0_inst_seg7_display_oseg7                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG7 -> system_0_inst_seg7_display_bfm:sig_oSEG7
	signal system_0_inst_seg7_display_oseg6                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG6 -> system_0_inst_seg7_display_bfm:sig_oSEG6
	signal system_0_inst_seg7_display_oseg0                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG0 -> system_0_inst_seg7_display_bfm:sig_oSEG0
	signal system_0_inst_seg7_display_oseg1                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG1 -> system_0_inst_seg7_display_bfm:sig_oSEG1
	signal system_0_inst_seg7_display_oseg2                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG2 -> system_0_inst_seg7_display_bfm:sig_oSEG2
	signal system_0_inst_seg7_display_oseg3                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG3 -> system_0_inst_seg7_display_bfm:sig_oSEG3
	signal system_0_inst_seg7_display_oseg4                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG4 -> system_0_inst_seg7_display_bfm:sig_oSEG4
	signal system_0_inst_seg7_display_oseg5                                                : std_logic_vector(6 downto 0);  -- system_0_inst:seg7_display_oSEG5 -> system_0_inst_seg7_display_bfm:sig_oSEG5
	signal system_0_inst_sdram_0_wire_cs_n                                                 : std_logic;                     -- system_0_inst:zs_cs_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cs_n
	signal system_0_inst_sdram_0_wire_ba                                                   : std_logic_vector(1 downto 0);  -- system_0_inst:zs_ba_from_the_sdram_0 -> sdram_0_my_partner:zs_ba
	signal system_0_inst_sdram_0_wire_dqm                                                  : std_logic_vector(1 downto 0);  -- system_0_inst:zs_dqm_from_the_sdram_0 -> sdram_0_my_partner:zs_dqm
	signal system_0_inst_sdram_0_wire_cke                                                  : std_logic;                     -- system_0_inst:zs_cke_from_the_sdram_0 -> sdram_0_my_partner:zs_cke
	signal system_0_inst_sdram_0_wire_addr                                                 : std_logic_vector(11 downto 0); -- system_0_inst:zs_addr_from_the_sdram_0 -> sdram_0_my_partner:zs_addr
	signal system_0_inst_sdram_0_wire_we_n                                                 : std_logic;                     -- system_0_inst:zs_we_n_from_the_sdram_0 -> sdram_0_my_partner:zs_we_n
	signal system_0_inst_sdram_0_wire_ras_n                                                : std_logic;                     -- system_0_inst:zs_ras_n_from_the_sdram_0 -> sdram_0_my_partner:zs_ras_n
	signal system_0_inst_sdram_0_wire_cas_n                                                : std_logic;                     -- system_0_inst:zs_cas_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cas_n
	signal sdram_0_my_partner_conduit_dq                                                   : std_logic_vector(15 downto 0); -- [] -> [sdram_0_my_partner:zs_dq, system_0_inst:zs_dq_to_and_from_the_sdram_0]
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0        : std_logic_vector(0 downto 0);  -- system_0_inst:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_write_n_to_the_cfi_flash_0
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0       : std_logic_vector(0 downto 0);  -- system_0_inst:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_select_n_to_the_cfi_flash_0
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address        : std_logic_vector(21 downto 0); -- system_0_inst:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_address
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn          : std_logic_vector(0 downto 0);  -- system_0_inst:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_readn
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data           : std_logic_vector(7 downto 0);  -- [] -> [system_0_inst:tri_state_bridge_0_data, tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_data]
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0       : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_write_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0      : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_select_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address       : std_logic_vector(21 downto 0); -- tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_address -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_address
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data          : std_logic_vector(7 downto 0);  -- [] -> [tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_data, tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_data]
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn         : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_readn -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_readn
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out      : std_logic_vector(21 downto 0); -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_address_out -> cfi_flash_0_external_mem_bfm:cdt_address
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_chipselect_n_out -> cfi_flash_0_external_mem_bfm:cdt_chipselect
	signal cfi_flash_0_external_mem_bfm_conduit_tcm_data_out                               : std_logic_vector(7 downto 0);  -- [] -> [cfi_flash_0_external_mem_bfm:cdt_data_io, tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_data_out]
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out      : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_write_n_out -> cfi_flash_0_external_mem_bfm:cdt_write
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out       : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_read_n_out -> cfi_flash_0_external_mem_bfm:cdt_read

begin

	system_0_inst : component system_0
		port map (
			clk_50                               => system_0_inst_clk_50_clk_in_bfm_clk_clk,                                   --                   clk_50_clk_in.clk
			bidir_port_to_and_from_the_SD_DAT    => system_0_inst_sd_dat_external_connection_export,                           --      SD_DAT_external_connection.export
			out_port_from_the_led_red            => system_0_inst_led_red_external_connection_export,                          --     led_red_external_connection.export
			zs_addr_from_the_sdram_0             => system_0_inst_sdram_0_wire_addr,                                           --                    sdram_0_wire.addr
			zs_ba_from_the_sdram_0               => system_0_inst_sdram_0_wire_ba,                                             --                                .ba
			zs_cas_n_from_the_sdram_0            => system_0_inst_sdram_0_wire_cas_n,                                          --                                .cas_n
			zs_cke_from_the_sdram_0              => system_0_inst_sdram_0_wire_cke,                                            --                                .cke
			zs_cs_n_from_the_sdram_0             => system_0_inst_sdram_0_wire_cs_n,                                           --                                .cs_n
			zs_dq_to_and_from_the_sdram_0        => sdram_0_my_partner_conduit_dq,                                             --                                .dq
			zs_dqm_from_the_sdram_0              => system_0_inst_sdram_0_wire_dqm,                                            --                                .dqm
			zs_ras_n_from_the_sdram_0            => system_0_inst_sdram_0_wire_ras_n,                                          --                                .ras_n
			zs_we_n_from_the_sdram_0             => system_0_inst_sdram_0_wire_we_n,                                           --                                .we_n
			tri_state_bridge_0_data              => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,     -- tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
			tri_state_bridge_0_readn             => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,    --                                .tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0           => system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,  --                                .write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address           => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,  --                                .tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0          => system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0, --                                .select_n_to_the_cfi_flash_0
			reset_n                              => system_0_inst_merged_resets_in_reset_bfm_reset_reset,                      --          merged_resets_in_reset.reset_n
			bidir_port_to_and_from_the_SD_CMD    => system_0_inst_sd_cmd_external_connection_export,                           --      SD_CMD_external_connection.export
			in_port_to_the_button_pio            => system_0_inst_button_pio_external_connection_bfm_conduit_export,           --  button_pio_external_connection.export
			USB_DATA_to_and_from_the_ISP1362     => system_0_inst_isp1362_conduit_end_data,                                    --             ISP1362_conduit_end.DATA
			USB_ADDR_from_the_ISP1362            => system_0_inst_isp1362_conduit_end_addr,                                    --                                .ADDR
			USB_RD_N_from_the_ISP1362            => system_0_inst_isp1362_conduit_end_rd_n,                                    --                                .RD_N
			USB_WR_N_from_the_ISP1362            => system_0_inst_isp1362_conduit_end_wr_n,                                    --                                .WR_N
			USB_CS_N_from_the_ISP1362            => system_0_inst_isp1362_conduit_end_cs_n,                                    --                                .CS_N
			USB_RST_N_from_the_ISP1362           => system_0_inst_isp1362_conduit_end_rst_n,                                   --                                .RST_N
			USB_INT0_to_the_ISP1362              => system_0_inst_isp1362_conduit_end_bfm_conduit_int0,                        --                                .INT0
			USB_INT1_to_the_ISP1362              => system_0_inst_isp1362_conduit_end_bfm_conduit_int1,                        --                                .INT1
			out_port_from_the_SD_CLK             => system_0_inst_sd_clk_external_connection_export,                           --      SD_CLK_external_connection.export
			out_port_from_the_led_green          => system_0_inst_led_green_external_connection_export,                        --   led_green_external_connection.export
			in_port_to_the_switch_pio            => system_0_inst_switch_pio_external_connection_bfm_conduit_export,           --  switch_pio_external_connection.export
			LCD_RS_from_the_lcd_16207_0          => system_0_inst_lcd_16207_0_external_rs,                                     --            lcd_16207_0_external.RS
			LCD_RW_from_the_lcd_16207_0          => system_0_inst_lcd_16207_0_external_rw,                                     --                                .RW
			LCD_data_to_and_from_the_lcd_16207_0 => system_0_inst_lcd_16207_0_external_data,                                   --                                .data
			LCD_E_from_the_lcd_16207_0           => system_0_inst_lcd_16207_0_external_e,                                      --                                .E
			rxd_to_the_uart_0                    => system_0_inst_uart_0_external_connection_bfm_conduit_rxd,                  --      uart_0_external_connection.rxd
			txd_from_the_uart_0                  => system_0_inst_uart_0_external_connection_txd,                              --                                .txd
			audio_0_oAUD_DATA                    => system_0_inst_audio_0_oaud_data,                                           --                         audio_0.oAUD_DATA
			audio_0_oAUD_LRCK                    => system_0_inst_audio_0_oaud_lrck,                                           --                                .oAUD_LRCK
			audio_0_oAUD_BCK                     => system_0_inst_audio_0_oaud_bck,                                            --                                .oAUD_BCK
			audio_0_oAUD_XCK                     => system_0_inst_audio_0_oaud_xck,                                            --                                .oAUD_XCK
			audio_0_iCLK_18_4                    => system_0_inst_audio_0_bfm_conduit_iclk_18_4,                               --                                .iCLK_18_4
			vga_0_VGA_R                          => system_0_inst_vga_0_vga_r,                                                 --                           vga_0.VGA_R
			vga_0_VGA_G                          => system_0_inst_vga_0_vga_g,                                                 --                                .VGA_G
			vga_0_VGA_B                          => system_0_inst_vga_0_vga_b,                                                 --                                .VGA_B
			vga_0_VGA_HS                         => system_0_inst_vga_0_vga_hs,                                                --                                .VGA_HS
			vga_0_VGA_VS                         => system_0_inst_vga_0_vga_vs,                                                --                                .VGA_VS
			vga_0_VGA_SYNC                       => system_0_inst_vga_0_vga_sync,                                              --                                .VGA_SYNC
			vga_0_VGA_BLANK                      => system_0_inst_vga_0_vga_blank,                                             --                                .VGA_BLANK
			vga_0_VGA_CLK                        => system_0_inst_vga_0_vga_clk,                                               --                                .VGA_CLK
			vga_0_iCLK_25                        => system_0_inst_vga_0_bfm_conduit_iclk_25,                                   --                                .iCLK_25
			dm9000a_iOSC_50                      => system_0_inst_dm9000a_bfm_conduit_iosc_50,                                 --                         dm9000a.iOSC_50
			dm9000a_ENET_DATA                    => system_0_inst_dm9000a_enet_data,                                           --                                .ENET_DATA
			dm9000a_ENET_CMD                     => system_0_inst_dm9000a_enet_cmd,                                            --                                .ENET_CMD
			dm9000a_ENET_RD_N                    => system_0_inst_dm9000a_enet_rd_n,                                           --                                .ENET_RD_N
			dm9000a_ENET_WR_N                    => system_0_inst_dm9000a_enet_wr_n,                                           --                                .ENET_WR_N
			dm9000a_ENET_CS_N                    => system_0_inst_dm9000a_enet_cs_n,                                           --                                .ENET_CS_N
			dm9000a_ENET_RST_N                   => system_0_inst_dm9000a_enet_rst_n,                                          --                                .ENET_RST_N
			dm9000a_ENET_CLK                     => system_0_inst_dm9000a_enet_clk,                                            --                                .ENET_CLK
			dm9000a_ENET_INT                     => system_0_inst_dm9000a_bfm_conduit_enet_int,                                --                                .ENET_INT
			seg7_display_oSEG0                   => system_0_inst_seg7_display_oseg0,                                          --                    seg7_display.oSEG0
			seg7_display_oSEG1                   => system_0_inst_seg7_display_oseg1,                                          --                                .oSEG1
			seg7_display_oSEG2                   => system_0_inst_seg7_display_oseg2,                                          --                                .oSEG2
			seg7_display_oSEG3                   => system_0_inst_seg7_display_oseg3,                                          --                                .oSEG3
			seg7_display_oSEG4                   => system_0_inst_seg7_display_oseg4,                                          --                                .oSEG4
			seg7_display_oSEG5                   => system_0_inst_seg7_display_oseg5,                                          --                                .oSEG5
			seg7_display_oSEG6                   => system_0_inst_seg7_display_oseg6,                                          --                                .oSEG6
			seg7_display_oSEG7                   => system_0_inst_seg7_display_oseg7                                           --                                .oSEG7
		);

	system_0_inst_clk_50_clk_in_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => system_0_inst_clk_50_clk_in_bfm_clk_clk  -- clk.clk
		);

	system_0_inst_merged_resets_in_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => system_0_inst_merged_resets_in_reset_bfm_reset_reset, -- reset.reset_n
			clk   => system_0_inst_clk_50_clk_in_bfm_clk_clk               --   clk.clk
		);

	system_0_inst_sd_dat_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => system_0_inst_sd_dat_external_connection_export  -- conduit.export
		);

	system_0_inst_led_red_external_connection_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => system_0_inst_led_red_external_connection_export  -- conduit.export
		);

	system_0_inst_sd_cmd_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => system_0_inst_sd_cmd_external_connection_export  -- conduit.export
		);

	system_0_inst_button_pio_external_connection_bfm : component altera_conduit_bfm_0003
		port map (
			sig_export => system_0_inst_button_pio_external_connection_bfm_conduit_export  -- conduit.export
		);

	system_0_inst_isp1362_conduit_end_bfm : component altera_conduit_bfm_0004
		port map (
			sig_DATA  => system_0_inst_isp1362_conduit_end_data,             -- conduit.DATA
			sig_ADDR  => system_0_inst_isp1362_conduit_end_addr,             --        .ADDR
			sig_RD_N  => system_0_inst_isp1362_conduit_end_rd_n,             --        .RD_N
			sig_WR_N  => system_0_inst_isp1362_conduit_end_wr_n,             --        .WR_N
			sig_CS_N  => system_0_inst_isp1362_conduit_end_cs_n,             --        .CS_N
			sig_RST_N => system_0_inst_isp1362_conduit_end_rst_n,            --        .RST_N
			sig_INT0  => system_0_inst_isp1362_conduit_end_bfm_conduit_int0, --        .INT0
			sig_INT1  => system_0_inst_isp1362_conduit_end_bfm_conduit_int1  --        .INT1
		);

	system_0_inst_sd_clk_external_connection_bfm : component altera_conduit_bfm_0005
		port map (
			sig_export => system_0_inst_sd_clk_external_connection_export  -- conduit.export
		);

	system_0_inst_led_green_external_connection_bfm : component altera_conduit_bfm_0006
		port map (
			sig_export => system_0_inst_led_green_external_connection_export  -- conduit.export
		);

	system_0_inst_switch_pio_external_connection_bfm : component altera_conduit_bfm_0007
		port map (
			sig_export => system_0_inst_switch_pio_external_connection_bfm_conduit_export  -- conduit.export
		);

	system_0_inst_lcd_16207_0_external_bfm : component altera_conduit_bfm_0008
		port map (
			sig_RS   => system_0_inst_lcd_16207_0_external_rs,   -- conduit.RS
			sig_RW   => system_0_inst_lcd_16207_0_external_rw,   --        .RW
			sig_data => system_0_inst_lcd_16207_0_external_data, --        .data
			sig_E    => system_0_inst_lcd_16207_0_external_e     --        .E
		);

	system_0_inst_uart_0_external_connection_bfm : component altera_conduit_bfm_0009
		port map (
			sig_rxd => system_0_inst_uart_0_external_connection_bfm_conduit_rxd, -- conduit.rxd
			sig_txd => system_0_inst_uart_0_external_connection_txd              --        .txd
		);

	system_0_inst_audio_0_bfm : component altera_conduit_bfm_0010
		port map (
			sig_oAUD_DATA => system_0_inst_audio_0_oaud_data,             -- conduit.oAUD_DATA
			sig_oAUD_LRCK => system_0_inst_audio_0_oaud_lrck,             --        .oAUD_LRCK
			sig_oAUD_BCK  => system_0_inst_audio_0_oaud_bck,              --        .oAUD_BCK
			sig_oAUD_XCK  => system_0_inst_audio_0_oaud_xck,              --        .oAUD_XCK
			sig_iCLK_18_4 => system_0_inst_audio_0_bfm_conduit_iclk_18_4  --        .iCLK_18_4
		);

	system_0_inst_vga_0_bfm : component altera_conduit_bfm_0011
		port map (
			sig_VGA_R     => system_0_inst_vga_0_vga_r,               -- conduit.VGA_R
			sig_VGA_G     => system_0_inst_vga_0_vga_g,               --        .VGA_G
			sig_VGA_B     => system_0_inst_vga_0_vga_b,               --        .VGA_B
			sig_VGA_HS    => system_0_inst_vga_0_vga_hs,              --        .VGA_HS
			sig_VGA_VS    => system_0_inst_vga_0_vga_vs,              --        .VGA_VS
			sig_VGA_SYNC  => system_0_inst_vga_0_vga_sync,            --        .VGA_SYNC
			sig_VGA_BLANK => system_0_inst_vga_0_vga_blank,           --        .VGA_BLANK
			sig_VGA_CLK   => system_0_inst_vga_0_vga_clk,             --        .VGA_CLK
			sig_iCLK_25   => system_0_inst_vga_0_bfm_conduit_iclk_25  --        .iCLK_25
		);

	system_0_inst_dm9000a_bfm : component altera_conduit_bfm_0012
		port map (
			sig_iOSC_50    => system_0_inst_dm9000a_bfm_conduit_iosc_50,  -- conduit.iOSC_50
			sig_ENET_DATA  => system_0_inst_dm9000a_enet_data,            --        .ENET_DATA
			sig_ENET_CMD   => system_0_inst_dm9000a_enet_cmd,             --        .ENET_CMD
			sig_ENET_RD_N  => system_0_inst_dm9000a_enet_rd_n,            --        .ENET_RD_N
			sig_ENET_WR_N  => system_0_inst_dm9000a_enet_wr_n,            --        .ENET_WR_N
			sig_ENET_CS_N  => system_0_inst_dm9000a_enet_cs_n,            --        .ENET_CS_N
			sig_ENET_RST_N => system_0_inst_dm9000a_enet_rst_n,           --        .ENET_RST_N
			sig_ENET_CLK   => system_0_inst_dm9000a_enet_clk,             --        .ENET_CLK
			sig_ENET_INT   => system_0_inst_dm9000a_bfm_conduit_enet_int  --        .ENET_INT
		);

	system_0_inst_seg7_display_bfm : component altera_conduit_bfm_0013
		port map (
			sig_oSEG0 => system_0_inst_seg7_display_oseg0, -- conduit.oSEG0
			sig_oSEG1 => system_0_inst_seg7_display_oseg1, --        .oSEG1
			sig_oSEG2 => system_0_inst_seg7_display_oseg2, --        .oSEG2
			sig_oSEG3 => system_0_inst_seg7_display_oseg3, --        .oSEG3
			sig_oSEG4 => system_0_inst_seg7_display_oseg4, --        .oSEG4
			sig_oSEG5 => system_0_inst_seg7_display_oseg5, --        .oSEG5
			sig_oSEG6 => system_0_inst_seg7_display_oseg6, --        .oSEG6
			sig_oSEG7 => system_0_inst_seg7_display_oseg7  --        .oSEG7
		);

	sdram_0_my_partner : component altera_sdram_partner_module
		port map (
			clk      => system_0_inst_clk_50_clk_in_bfm_clk_clk, --     clk.clk
			zs_dq    => sdram_0_my_partner_conduit_dq,           -- conduit.dq
			zs_addr  => system_0_inst_sdram_0_wire_addr,         --        .addr
			zs_ba    => system_0_inst_sdram_0_wire_ba,           --        .ba
			zs_cas_n => system_0_inst_sdram_0_wire_cas_n,        --        .cas_n
			zs_cke   => system_0_inst_sdram_0_wire_cke,          --        .cke
			zs_cs_n  => system_0_inst_sdram_0_wire_cs_n,         --        .cs_n
			zs_dqm   => system_0_inst_sdram_0_wire_dqm,          --        .dqm
			zs_ras_n => system_0_inst_sdram_0_wire_ras_n,        --        .ras_n
			zs_we_n  => system_0_inst_sdram_0_wire_we_n          --        .we_n
		);

	tri_state_bridge_0_bridge_0_tcb_translator : component altera_tristate_conduit_bridge_translator
		port map (
			in_tri_state_bridge_0_data     => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,      --  in.tri_state_bridge_0_data
			in_tri_state_bridge_0_readn    => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,     --    .tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0  => system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,   --    .write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_address  => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,   --    .tri_state_bridge_0_address
			in_select_n_to_the_cfi_flash_0 => system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0,  --    .select_n_to_the_cfi_flash_0
			tri_state_bridge_0_data        => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data,     -- out.tri_state_bridge_0_data
			tri_state_bridge_0_readn       => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn,    --    .tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0     => tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0,  --    .write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address     => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address,  --    .tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0    => tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0  --    .select_n_to_the_cfi_flash_0
		);

	tri_state_bridge_0_pinsharer_0_pin_divider : component altera_conduit_pin_divider
		port map (
			in_tri_state_bridge_0_address    => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address,       --              in.tri_state_bridge_0_address
			in_tri_state_bridge_0_readn      => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn,         --                .tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0    => tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0,       --                .write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_data       => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data,          --                .tri_state_bridge_0_data
			in_select_n_to_the_cfi_flash_0   => tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0,      --                .select_n_to_the_cfi_flash_0
			cfi_flash_0_tcm_address_out      => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out,      -- cfi_flash_0_tcm.tcm_address_out
			cfi_flash_0_tcm_read_n_out       => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out,       --                .tcm_read_n_out
			cfi_flash_0_tcm_write_n_out      => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out,      --                .tcm_write_n_out
			cfi_flash_0_tcm_data_out         => cfi_flash_0_external_mem_bfm_conduit_tcm_data_out,                               --                .tcm_data_out
			cfi_flash_0_tcm_chipselect_n_out => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out  --                .tcm_chipselect_n_out
		);

	cfi_flash_0_external_mem_bfm : component altera_external_memory_bfm_vhdl
		generic map (
			USE_CHIPSELECT           => 1,
			USE_WRITE                => 1,
			USE_READ                 => 1,
			USE_OUTPUTENABLE         => 0,
			USE_BEGINTRANSFER        => 0,
			ACTIVE_LOW_BYTEENABLE    => 0,
			ACTIVE_LOW_CHIPSELECT    => 1,
			ACTIVE_LOW_WRITE         => 1,
			ACTIVE_LOW_READ          => 1,
			ACTIVE_LOW_OUTPUTENABLE  => 0,
			ACTIVE_LOW_BEGINTRANSFER => 0,
			ACTIVE_LOW_RESET         => 0,
			CDT_ADDRESS_W            => 22,
			CDT_SYMBOL_W             => 8,
			CDT_NUMSYMBOLS           => 1,
			INIT_FILE                => "altera_external_memory_bfm.hex",
			CDT_READ_LATENCY         => 0,
			VHDL_ID                  => 0
		)
		port map (
			clk               => system_0_inst_clk_50_clk_in_bfm_clk_clk,                                            --     clk.clk
			cdt_write         => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out(0),      -- conduit.tcm_write_n_out
			cdt_read          => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out(0),       --        .tcm_read_n_out
			cdt_chipselect    => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out(0), --        .tcm_chipselect_n_out
			cdt_address       => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out,         --        .tcm_address_out
			cdt_data_io       => cfi_flash_0_external_mem_bfm_conduit_tcm_data_out,                                  --        .tcm_data_out
			cdt_outputenable  => '0',                                                                                -- (terminated)
			cdt_begintransfer => '0',                                                                                -- (terminated)
			cdt_byteenable    => "1",                                                                                -- (terminated)
			cdt_reset         => '0'                                                                                 -- (terminated)
		);

end architecture rtl; -- of system_0_tb
