`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eu0A6FN1D763eFAO04lO75wSh+q2FJ09LrYcDlK3ukdWb822zd/YORjkOQ8eLBJg
/+Clg9QlAGoN9AQYDS65AQPR2GnuU3QHqvaKbIfyC8BOnUXLwYk1IeAg6frgc3gc
oWQzD4yj4BHqTXY1uMo5KeJUckRg6yimjMjyvWF6QzEVgJNcqFhbmdc5FjbwSeck
vuv2mzC1E2mEdRq30kk3oOm1QYopjPL3wt2zf1vHX6U=
`protect END_PROTECTED
