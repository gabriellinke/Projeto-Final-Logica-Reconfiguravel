`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJY/oQ+Y+sog4ZEeqX5oOFzzhtpGGO78sTBz6rPoF/94N4bH+7yNc6fnEywNBazt
6lgHb9HfiUev5TWKWd19nXdTcAjbockSbknkRvngRMfBjhySMn/HLk00PrAERar/
yu8fUUADOJ3k9AnhZ+t8H1/gvvW8YBpP02sj2P4uS8SIiONUzZ/kkedPlOHSuEJY
z5MJ45aRaST259zp8aGJqH7jPS4c0MjmiZVFy8GHktJ8JLtdTVtVOK4GrGQxUEMU
ggPk1xwUEdpjujk7qw6SXcJ2AoPSgFsux0e+SFhm3Ct4GhUgkqKgJBNL+Wkap1gd
1XcLWZRQKsIOoO2aX4mDwASU6inX5LRGinZHl/2cPmUAhBpNWPxyj/ew3U8fPyw2
aS1/DdPn2V9d6d2FQ/TIzLiMdcFfSi3oVlN2dS03Y+R6phn3u7rNUT3UPOGV95kJ
eMgvrMUscCFLLcs9SxCUkzQGJLf9L40gwdeTBinpLpqtBZJtqfopQC9ZgDSaxwe6
VVjs2jfxn7TtjgiNy7rQuG2KR5aFOCTbBIrmpFcrUYE8YNHWNDsBXs00hHFrCMGZ
PbYN3NPRc/opbPBiFluk5HTLzojPIJi74LOXT/SwEl3uTuPd60CQ1yzJIFxyVEx1
YWCjg39F9qQ4XRvYzIWTp/p8ipCp+hlsBDTg1kTzFuI7aiLqPk08R57kudrAXwGu
U89hylgd+KlUNJ+3U+OP0KmCSV1OynttYEH513vK1Xel/VEKI52HqY11QGnr9QC8
ZYJNTYYFItZbcpLl/nhQBgjRU0V0678VcTyXQvPK3AHj1KgDdRUxn2OzGmBnvpvb
j4uPvFjDqcG3BzW96dwgcM39j5laR8yTJnA6xx8EJ1idMHEv+tPfIa9riCHTT+mN
mCvHnEfus/x7cWqiweGf8f5SRgOrfSUabG6+rAlAJ3SF5uqUxNA8TvMgnRkb0ubq
8ku0xKLUXCuqT3EcXTuHmnY0JDwxB3XXx3oJGUynv0Boi2EpRFuQGd113F2FXSLf
SerlxPOBXtsESAwYbeyCshPap8JE7Ic0r6/xi0QjODPPfCYkop3WLa5K/KYaG7tZ
flTxI3n/G8t4df6vilG/V3D2hbazGCE3EsbKV6y0n5xgeMzNO67vVPNUwcrNFnXW
0qzCV37g9vph43uZHBlO0KuHkufqhXwHShzvXgE7BnSqwG5z9NKnlHSYzLz0xd4Q
bfCvhBjeLItlvuy00CV+19Vj8gB7QQUBtBg5nOwNmLntpK5/Sr4Bul0k99Vfbz9H
eT1tOJat70f2aNfEe0YtrrAHGW23qkJ180Unq2TmYw/fmn1lvISSG1yh3o768Vd3
09PxfWX4sQTKC+N3PyGop1W6U7ZpfyI/G5xgy56tcSb/y0R8Sy/YJjFcb0p9JHil
MCjOodOnxK34Wn6O9ijqv0KwEIBLWe02YwrOV2dxzjqyzL/TIzekV45+afVmtAT9
Nmie+GpHzyfuKF4ngb8F4PX6JNRFTMAMIyEVRVEOUT/Dty6HYF+YGjl7lysNmIj+
1+HosI9YoUuR+JzqI4A/WnyH0nQ8eCUbTj/sXkf8KtrcXdZzkGT4NLceMPn3juah
RHNB5srBbRzZ6Q01cmUAOUqu/4bPiDlOKDhf6c30Lhk2dLh8kjJdzxNJY99dXn0O
ZrrqPuxNqY31v5KnRbfxB15y+rr1T380PsRW60L6GidZlM/VVy3cy3/w8o1BQJma
b8UuhHfVUUThYh2gaQcjcg3+SHFH777G2QWMR1x0Ysop9fha0mOtP4sMzkVhjMW0
Ac/+QEa21jeU0VgWuvLL5USUH/0CbnKIFK+uHS6RNY0AP8FyPc+e65s8ZynBfSHu
STLLTF2LqK7r3RS2iwuqG1aZ+1RjvqQPXrHg6olet1DfhhYFq8Cb/0Qly85+lj7/
bbEMsXLuSxoXP77juKbYGuKlYgT7BAzOlfRmu2DjHO+3ILr9uSlTeA5L2pvuLZWW
iH6l5jIDYq7WaPwS0YOluzeqF57ojUND2TExVf1OfVt02LXRn1GpPE4hZAMPVVRX
HyVEnb/un1S4etPk0iC5Tq1eHP+DzB7RZ8YheaWSXoZFA2eDxzNAnB+t34y96mzk
VPdhuOORCoetzQMG80licPLWR0s6fnft0C6717kbDb5vdR5nUIo5c0Uw5QWDdzuQ
04NjeC1EdWsBxH41S1wbBCQvBku7Nkl8a85ihFr/97EtWgfFVo3WeGVc/YizvFzL
C/4tc9cXkz01zGWxC/67eElz1G9/GQ3gvOb4gIggrrDDaili4YnGgBuEa+kFevHD
TEQ5Ayk4i212SAmj448ufbOP/tbN4LFAJnOIUy/NB9M4kRlhMNt418CyFsq2e80W
c7JZCiA2ZqmfsAJzQOUGDFVqQiMhglH3upOjN71ngmitjjnNMs3bSWWcTzb5o5sT
dSyMWyeY6d8ivz0/J80RBxfbB/1XrA54/gNUiMcarn+M4tSKf8XXy6mWOB7Qzq/4
ksd4Q/ljAKHrDnj4lJLfdDRj8uQE3QllC8MpY9exnKcEoz2dt9NZWRVTC0rfZjWu
GyK7AhEHkKYPvbDJ14DXwnrqAA+flRWEyiomjTOCEatG2whxOTkYinicSD2Tf/3p
Qe7bkIG7w4Sr6Z1Q3G7GM9EnN2CU8D9ZbP+dmlJluH97Dt7nMbc6FQQ/Ta+sA6l0
vdcBBWplAKKg16RQOSJCaQqqjSOsnzinWhTQmYYls0FDDtQiYPOZk1vF7fb8gTjZ
Vif3MbKKELSteUo98mvZProczeV2ljObSm+6Z/PpUpp+NsR7eM+C6JcBTgpXo5Td
Y6XVpVitJNiVMDp2Pe34CKIf1L+s+xtrdg84uz6j6DmhWqpqwq3ozF9UpCYz2qPX
OTL9kIVf0LxPSoY1EBHrlETy+m6p2I/r21mAAPtQYXBvwv3C7fW4VyZTekHnPrNL
57YR1JVsh6md6TnpN7DBmx7XD7XZsOh7nQSFxgqPQzmJN//aylzXRj4fAVnpO/L3
wxrSECblejYPWyjdtMmpXuKDwSqjv9HE13uELnMRUs8P68qenI0+3ZBv8wNx00aR
Z6yzBEmYxp2K6WuBAE6L0byeTA28TbPkbUsFWp/YCHh3Q/LR/IH4pbAGPs3ysnzr
XSFW6BtzBNa+AWKWzVvnWOCbgdoqQ01DKLUo2FPbMTuj2NsKpvyBZt4sf99PJ2io
FgPxdwPDuS+WknSEBWIbeg9kuQhKnPYfgVNdut6rZlYFGs296N75aqJLGF9ZXsPF
O8IDAFZNd8Wpa82Zn6tHqnc/BirYmkwDkEfb7eZ48h9AkEkFj0pgzzeDXOXDgr5G
1Foh/ZRkkmeHp7j0eMfs+U/zZTaNNFbndnIrQZHQ+jUagh1pFZxR7iknSUlNW9mr
ZHGdKikk2UbcGs/PaKvSJ2PuRG9qJ5WM9mJQikbEzd+ULWKl7BsR0lmaiFO3PHcf
9yTamrGDSYCGI1Eg7Gqu3Xho8YaHEvgRxZ2jzNq89SlbAFXzYScdh3maz/erpYz2
re7jxovGVF3mMBdfA13SWgDkjwbzbJjlsO6s+tSr10MUFatIOp9htEKcrZAsM8BA
tpI+Z8z9op6y8rf/Y3toxYLlaPToFdDihl8Xflfyy0xrz3EWcnB3/tmddQzWo1Nz
AMjBbbQmugY1xL4yZBWRKPAgNr3n5fezuYnc7BBvgyZZfAaQO064DeJGvS0rtoDw
wAVsL5EpIxKOVjWjSsiDJS6l5G2f8/k29a5GRr7uZAAHY+aWZuSz73mfwcTTexwI
li6JvnSBWayMIZap0PMgBkYm/2EhQfcu2Z9ZTUK9C619AAZ7OpIzRY35ttoZtysT
n/fh6dXONwLd59Uc0RrsSH2WNa93P5HXxD/r1+yLD7Xf98Y1Nv46qj0Oqx47v2SA
dxNOVmuvQ8K8UU/H+db+jEojlRt2TE8jp4uvAGSb7+D6HE2v1guzA/NABlmuWPoz
eVWS4ZONq1JBBJG6wYSMVMZ8gJt6P91SdqzeTWRniJz9LvMeuawupbkZDLupdK4T
ABmEbmeIzPm42L0a8lCypL7gGuwhOl57yg9t8doiqcbcsJXsd+2Wv0p3M7ObFdh+
krlSUSwIbcyRi/rvo7UrSieyCJUI0lgorGHQAdJJWxF0mTqStipRzSJuKNf0E274
+4BGQZYtHzgUEjlPfdb9WqrD/H3yE/+CJ0ETBryZyCCOmHz9Wc4Y749+lg5HLsZY
2bDR/IGGBTADBRO/0J1pHX1CvnKIFXyCo20pBeNdUz+uutxVoPHeyRGZtV2mmQyu
FUVrGZxIur/6a3oql9aW5Ld8dRn2qSwhyyAmN/5HEtaen/TicdGihQmV1CHjCmRG
VPhmIM4Fo88v1wg56CML6HI6aUlgEvjdiiN9m+UNO9pKlQSOtYPUOOEY3u0RLr2F
dJO+bJBmuWqYxA9G6HhHJ6kqVEdbGfam7Fvapur4VZRAzptNFZk+aeoD/36ogeZJ
SVlakTeP7LK9L7+l4KlNOAgPw0ieh7U09yN9KGEKWM912RzMguS/RYxkiOXeRb9j
o9/t4VYKsslD4g5n0ldjF76NsySBKN87/MLbZVq2Cg+09jRoDOU9t9seK7HOfI0E
`protect END_PROTECTED
