`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/ouXLXQKLeRW7FhIg58sAKlmAXjTGhCQ8ABXTbuNIPTxlvSiU4OxCHrs+WbzxBK
ZPs4pFOsNdWPWUlITYNXwC9qr18ayvU/It/zIwl32A/3s0MyRUE3Z4nxpN81+Htf
1JXzhL7jZSpDSv/gDuv4/cv2ebfZFXk5sO7sjNsqe641nVVMSaJGGeV8gIyKFZNC
dc8lMN9kM6qoW+48OlGrsUXcY5YYD7p6YpIDDH8l1/DV8CxJt/eogM18XFaci2tF
Vf/iLVSgiI1cp5MwSstAuo1u81w2M1kbJHxkzB8e7UPpi1xJy1x7i7bzwF8LOX1a
stL/L/Tvz5Z2whDU5+Hvbb0qGuJv1786SU25ZpXGsHpnAzYw/iSZfdo+yhh8htY7
b5D9fPu9FPzI0BpIYukYKEh8HrZTEJ1urjjWibQ23SU6G1zZusrGijsTzKJZjPoP
HO60FFPb3b7KkPzv2hU17coNMfQk8aFXGrfJjVMndi6r8aYMj7moloF/IhyklExW
gMuvicVMLlouBWxILL+uQdveh68gOl3tz44kSFZYm9LhFR1lq8TsyCjNpoTacEQV
LWhq6oXBoKzjNTH7X40yA2bUZ/2O2vYdBpfcgfLFMN//fdcB1S8FBuoI+eJG8R2y
2dMd3dcgX3wNVJpBb8+n4MqroiHzQI+k/k7dKsfwIJ6D0ji/UXpG9+PW1w8DbwNh
z3qcGC0Q5sNUAM4JEq1zK+fW/Jf+G3Awi/NCqaNfdC38OhBaprqOO5LnM9dAJt3r
K+x2YFbxF0bS9acisN7VTrXtPtpyuc6/YNQ78kNfiarU3yoN5xk/R7ykAWxUJXNO
c5lOeOOadlsg59fhMO8MYsC12skXhvdKHKhb76Lu36miixckQNnnTfUqRA3pNcAx
U71ekkY6i4mUxrK+T9PvVFWZaIkWyD6U5HjdSSWsuO2r48nC8vdgStpb8+tjflgE
45TwxyIu0C+sxNq/n6erIreKTRZLa+vnpHEbzJXhLvC7Mxbfo6f4xYb/6YoMzBJ3
yyRikjIwSKpegGrJJa76s5XbcxvDZeUuwmtEX57kSX7TSierciOEoTSey+lF7pIi
k6Q6v+9SUi2UV5RW6g4FEvQk/emUHcHykfiHOQ9bwBJp0XSO0GhddCU5ODpwUlP6
bcuBpdpoXpleFzFZDUc/vikHrGMAsAs9hWnQge6WeTdSFPCPLXGQcbS33Gxd8zow
qCA4PSexg+aNvubFzCyCSNI3xMNJqJ5gvMOSBILKRvALla3LqQuSLWmXooM+Pj1p
UJ7iDigZQk2Nj6HMbFcmzGqpdy+X2Ve7y7fGSBp9YeF4ejG/ODfnTnuDgpqk0NXm
f+QiWfclOC8ktXzUl//PLB9vNd7C5BpjEHIBySsBJo4rQ+C1CKkhrAJqea0GZYvs
EweDtE1GG/CF/LEX4wMefKQqWsZ3u25DRr69SJ8lhywAMgx+STgXaFCodBnnU6sL
0Lfh8xm8PGBhcqw8VcYW65Fe/PrJR7ybDtWrzzLxz7GFNSUdLiEbpUEAZlsVBV5A
PVCDPp1iwd7sKLOeWeaajw0GXBVa2wtcl02QEiIK/yzPCRyUd20FEjtANUjOGqIB
Els6SkiQTuANDDSIaQIxV7JJdEcotXz3huFfSTpEmBoQtSI1toqrTknmdF5MYL8P
DSiFtXJ8gNOmqjcwbo6lTprh1RTuH4WIa0A9lECJ5qG4K4udhGVhlbfMHQDkaPYN
f5HTCHTis2bRVbQAgJaxowDeDo+oVTwnwzqTfNiK/byXnCvnOYHxqs55a6PhtR4x
5yic28JtnpPyQ84EHauWs8Pt8TTdXoujhtbSN4ZyJXSmg0JrDKiuJ9ptN90O5fzf
wwAGs4WAGl0gUql5qeAyiGiMQo1pSitV4sst8gZpJaJ5mLDe3CM4UgH/vkNKBENt
DrMa9qaWyPXUsQt0XZsD4UIeEa+w89XWhtJwOBKPjySIGmKSXRg1fthUChxXxsAH
YqtabUjtcKqN9RMEbHboiT6VOKRtl67l6vcmc5CfnwuMHYrWPM695IIYpFIPYmBn
L3eZQf33gKei9GI9eZgmFrI6ug3UDLb8pQKmWD1ZQMcuZZvFL25sxgU1bSc3GvkQ
78OVN+p3vY3PsKCSkLugpWTQ2IKfjuucbecNFBYRpJpsl2yv8VTsuTBn3JaFRQEG
vjwL7E5/2GUJgmYNBXOuXmYncgfq1xVr+xGzLuLLDZCGvp4QFH6dPosha49zJ6a+
lR8BXcWzxZF78wp3CAv/HbAG+v04aMdSLJrIwXlx/jr16MwhXLUJMYqyYkt8GVGL
VaJzOKWaLv8qTXWWssiZ2ooKpa4GSTIAYV1ztYkT4G7AEjVud6xLLXJ4F9P4mZGh
tskGcf+s4/L1kpMb5arQx/1fKaCD9e4uvRCCohO6imaiawacOUkMhWO2Nld4Si9C
Dz9Q4JfMPM19KMQCQTKDozQDdAlkemQK/hcHMEYkwTUN78guKmNTX8c1MUiaU7dd
iKx9Y/wvN8n1p4Vx8k63f7uBFp0jiAw7h5o7yZ6mD3cjdM/tGTLuxYz/Pr04/kNF
1fJ3rVCm8030LLntGF5I470E0u0DxBGhV3IphOuvyXuJh1pFxtPuZrIgUr+nM+Gc
wFG7iYxSaLr6i0EuWvqM90ZitUeIgLsnFopqWDWaoMQ+RykapJ0GRNGF0ZivBcgc
GqHmEcAkA0JGEQHEgr+73QFYpG2wDoCXhLeB6/6PPOeZ5eaI+YQf3U8wv137J+y4
VjaNzF+zWGZ+kKG0GtpVFgpDwdW9HZcJ+qDNIs+me1Z0OxovcK6qSR6fl/w6oV1V
Q11qWHmba2KrmthbHh3q8rx1tNSOHYjTQRqL4xc49d9K7T3nDxnKOltJ7G/ighS8
vhgecD32HrQm1GNTR5+T1Hl4ZNdJza7QBcUVzr/OCrrRYwBdqj07k6Hq7o1/CV2f
PWFNJGbuq5EgfAUd47BnJDYXCrkUhKG3otr5HHS/+dKcAlQiX/BuYJq6qfrs3F0I
YvpiLoU+CvbwP7QuVjF9+f9Y6WgltmMucBM31yB38Pp+qXEX9evwuXlpta4VgyEd
0+j3zFpuWCxK2DwzIfrDeyMdrT9YjIjtsaZM28hee14gAoewKaA5NXYp+06MZIlY
Yy4YYr/SR64uFamfz6GKCiRCtMt8gPvL1qR+4DdVW3mP9/2Vw2wPMpYzy3adgV1R
EkrSnaVX1wGjRR2SXKXqatvbqfrgA7Vuye4GLM/IqjgmL1QEeMdq/FfbqZ1NGIST
DD5RKaIn0ACz2M64Br10TZi67SHXvXEZokuiIjyVWEHU7K7Xb5nLNLoZVIKrjGM9
LxAThUq9LH+QCvmYRGDtYib5Zb7BEa8s6vkDZQ8/sVVeLnGb6c1DJjeVhpBBly0s
/HncSC4zMNmTH1hkvkDq3KtJzCPEnuZdJD3VJCk+HFB72TurxIfVsguE02SMMD+h
MiWwjNjQPnkXRPIZZQGez5bxrF/BMDmX9rmAdKJnPfXENPiY6YgoaSaGwOlpDwuk
KOAfNR4QUinHG3D+HGDri8UCSy0YSQ11C8SVfvwMTVR2GMsQPE4X6uwXfTvkhmxe
fPOQUK8hdeM9AYEJzeoWgdzsdqM2vTptQj/gd/F1acgSNjtCxOVbbOpKsAMCWRaJ
kYkTUw+6m2S7aublPkjLFg==
`protect END_PROTECTED
